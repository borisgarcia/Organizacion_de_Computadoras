`define ADD 6'h20
`define ADDU 6'h21
`define ADDI 6'h08
`define ADDIU 6'h09
`define SUB 6'h22
`define AND 6'h24
`define ANDI 6'hC
`define OR 6'h25
`define ORI 6'hD
`define SLT 6'h2A
`define LW 6'h23
`define SW 6'h2B
`define JUMP 6'h02
`define LUI 6'hF
`define LB 6'h20
`define LBU 6'h24
`define SB 6'h28
`define SH 6'h29
`define LH 6'h21
`define LHU 6'h25
`define BEQ 6'h04
`define BNE 6'h05
`define BGEZ 6'h1
`define BGTZ 6'h7
`define BLEZ 6'h6
`define BLTZ 6'h1
`define NOP 6'h0
`define SRL 6'h2
`define SLL 6'h0
`define SLLV 6'h4
`define SRLV 6'h6
`define SRA 6'h3
`define SRAV 6'h7
`define XOR 6'h26
`define SLTU 6'h2B
`define JR 6'h8
`define SUBU 6'h23
`define XORI 6'hE
`define SLTI 6'hA
`define SLTIU 6'hB
`define JAL 6'h3


